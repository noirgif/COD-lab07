`timescale 1ns / 1ps

module EXHU(
    output exc
    );
    
assign exc = 0;
endmodule
